module not1(y, a);

input a;
output y;
assign y =! a;

endmodule